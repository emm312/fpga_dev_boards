-- emacs 26